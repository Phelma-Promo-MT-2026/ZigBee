* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 10:07

.SUBCKT TOP
M$1 \$3 \$4 \$2 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
R$2 \$1 \$2 ptap1 A=0.6084p P=3.12u
.ENDS TOP
