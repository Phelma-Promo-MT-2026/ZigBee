** sch_path: /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/xschem/Zigbee/LVS/LAYOUT/test_capa/test_capa.sch
.subckt test_capa VIN VDD GND
*.PININFO VIN:B VDD:B GND:B
XC1 VIN net1 cap_cmim w=6.99e-6 l=6.99e-6 m=1
XM1 GND net1 VDD GND sg13_lv_nmos l=0.13u w=0.15u ng=1 m=1
.ends
