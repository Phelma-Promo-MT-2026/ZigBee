* Qucs 25.1.1  /home/userproj/microelectronics/ProjetZigbee/ZigBee/PLL/PLL_verilog_A/VCO_FDIV_test.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"
.SUBCKT VCO _net0 _net1 

NX1 _net0 0 _net1 vco1 
.MODEL vco1 VCO()
.ENDS
V1 vin 0 DC 0 PULSE( 0 1 0N 1N 1N 1M {(1M)+(1M)+(1N)+(1N)} )  AC 0
XSUB2 vin _net0 VCO

.control

tran 5.02513e-05 0.01 0 
write spice4qucs.tr1.plot v(vin)
destroy all
reset

exit
.endc
.END
