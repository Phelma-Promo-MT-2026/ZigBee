** sch_path: /home/userproj/microelectronics/projects/ZigBee/LVS/xschem/BGM_AA/NMOS_RESISTANCE/TOP.sch
.subckt TOP VIN GND VDD
*.PININFO VIN:I GND:B VDD:I
M1 VDD VIN net1 GND sg13_lv_nmos w=0.15u l=130n ng=1 m=1
XR1 GND net1 rsil w=10u l=10u m=1 b=0
.ends
