* Qucs 25.1.1  /home/userproj/microelectronics/projects/ZigBee/PLL/Pompe_Charge/Bascule_D.sch

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_pmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 
X1 d g s b  sg13_lv_pmos w={w} l={l} ng={ng} m={1} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout}
.ENDS
  

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  
.SUBCKT NAND _net3 _net1 _net2 

.LIB cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2

Xsg13_lv_pmos1 0  _net0 _net2 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos2 0  _net0 _net1 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 _net1 _net4 _net4 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net4 _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
.ENDS
.SUBCKT INV_2x _net1 _net2 
.LIB cornerMOSlv.lib mos_tt
V1 _net0 0 DC 1.2
Xsg13_lv_pmos1 0  _net0 _net2 _net1 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.6U l=0.13U ng=2 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net1 _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.ENDS
.SUBCKT NAND3 _net3 _net1 _net2 _net4 

.LIB cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2

Xsg13_lv_pmos2 0  _net0 _net1 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos1 0  _net0 _net2 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos3 0  _net0 _net4 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 _net1 _net5 _net5 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net5 _net2 _net6 _net6 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos3 0  _net6 _net4 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
.ENDS
.GLOBAL 0:G



XNAND2 _net3 _net4 _net5 NAND
XSUB5 _net6 _net2 INV_2x

XNAND3 _net7 _net8 _net4 NAND
XSUB3 _net9 _net4 _net1 _net8 NAND3
XSUB2 _net8 _net9 _net0 _net6 NAND3
XSUB4 _net4 _net7 _net1 _net6 NAND3

XSUB1 _net5 _net3 _net9 _net6 NAND3
.END
