* Qucs 25.1.1  /home/userproj/microelectronics/projects/ZigBee/LNA_grille_com/akrxm2a/SchemaCG_LNA_Single.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  
.LIB cornerMOSlv.lib mos_tt

V2 _net1 0 DC 1.2
Vin _net4 0 DC 1
L1 vout  _net5 3n
C1 _net5  vout 1.41p
R1 vout  _net5 500
Rs _net4  _net3 50
Lb 0  _net3 3.25n
Vdd _net5 0 DC 1.2

VId vout _net0 DC 0
VId1 _net2 _net6 DC 0
Xsg13_lv_nmos2 0  _net6 _net7 _net3 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=10U l=180N ng=5.88 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net0 _net1 _net2 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=10U l=180N ng=5.88 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
V1 _net7 0 DC 0.6

.control

op
print i(VId) i(VId1) v(vout)   > spice4qucs.dc1.ngspice.dc.print
destroy all
reset

exit
.endc
.END
