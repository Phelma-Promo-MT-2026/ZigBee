** sch_path: /home/userproj/microelectronics/projects/ZigBee/LVS/xschem/BGM_AA/NMOS_SIMPLE/TOP.sch
.subckt TOP VIN GND VDD
*.PININFO VIN:I GND:B VDD:I
M1 VDD VIN GND GND sg13_lv_nmos w=0.15u l=130n ng=1 m=1
.ends
