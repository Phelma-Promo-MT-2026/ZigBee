* Qucs 25.1.1  /home/userproj/microelectronics/projects/ZigBee/Techno/carac.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  

.LIB cornerRES.lib res_wcs

.LIB cornerMOSlv.lib mos_tt



Xsg13_lv_nmos1 0  Vds Vgs 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=10U l=0.140U ng={W/L} m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
V2 Vgs 0 DC 1
V1 Vds 0 DC 0.012926

.control

op
let Ids = -i(V1)
let gm = deriv(Ids)
let gm_sur_Ids = gm/Ids
let k = 29.4
let gm_sur_Ids_sur_k = gm_sur_Ids/k
print v(Vds) v(Vgs)  Ids gm gm_sur_Ids k gm_sur_Ids_sur_k > spice4qucs.dc1.ngspice.dc.print
destroy all
reset

dc v2 0 1 0.0126582
let Ids = -i(V1)
let gm = deriv(Ids)
let gm_sur_Ids = gm/Ids
let k = 29.4
let gm_sur_Ids_sur_k = gm_sur_Ids/k
write spice4qucs.vgs.plot v(Vds) v(Vgs) Ids gm gm_sur_Ids k gm_sur_Ids_sur_k
destroy all
reset

exit
.endc
.END
