* Extracted by KLayout with SG13G2 LVS runset on : 11/06/2025 11:49

.SUBCKT TOP
M$1 \$3 VIN VDD \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
R$2 GND \$3 rsil w=0.5u l=0.5u ps=0 b=0 m=1
.ENDS TOP
