* Qucs 25.1.1  /home/userproj/microelectronics/projects/ZigBee/PLL/PLL_ANALOG/PLL_ANALOG_Total.sch
.INCLUDE "/usr/share/qucs-s/xspice_cmlib/include/ngspice_mathfunc.inc"

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_pmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 
X1 d g s b  sg13_lv_pmos w={w} l={l} ng={ng} m={1} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout}
.ENDS
  
.SUBCKT INV _net1 _net2 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2
Xsg13_lv_nmos1 0  _net1 _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos1 0  _net0 _net2 _net1 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=2 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.ENDS
.SUBCKT NAND _net3 _net1 _net2 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2
Xsg13_lv_pmos1 0  _net0 _net2 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos2 0  _net0 _net1 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 _net1 _net4 _net4 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net4 _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.ENDS
.SUBCKT INV_2x _net1 _net2 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2
Xsg13_lv_pmos1 0  _net0 _net2 _net1 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.6U l=0.13U ng=2 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net1 _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.ENDS
.SUBCKT NAND3 _net3 _net1 _net2 _net4 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2
Xsg13_lv_pmos2 0  _net0 _net1 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos1 0  _net0 _net2 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos3 0  _net0 _net4 _net3 _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=0.3U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 _net1 _net5 _net5 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net5 _net2 _net6 _net6 IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos3 0  _net6 _net4 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=0.15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.ENDS
.SUBCKT Bascule_D _net3 _net2 _net0 _net1 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

XNAND2 _net3 _net4 _net5 NAND
XSUB5 _net6 _net2 INV_2x
XNAND3 _net7 _net8 _net4 NAND
XSUB3 _net9 _net4 _net1 _net8 NAND3
XSUB2 _net8 _net9 _net0 _net6 NAND3
XSUB4 _net4 _net7 _net1 _net6 NAND3
XSUB1 _net5 _net3 _net9 _net6 NAND3

.ENDS
.SUBCKT Diviseur_par_2_digital_symbole_ _net1 _net2 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt

XSUB3 _net0 _net1 INV
XSUB4 _net3 _net2 INV
XSUB2 _net2 0 _net4 _net0 Bascule_D
XSUB1 _net4 0 _net3 _net1 Bascule_D

.ENDS
.SUBCKT Diviseur_par_2_symbole _net3 H HBarre 

.LIB cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1.2
V2 _net1 0 DC 1.2
Xsg13_lv_pmos1 0  _net0 vin A _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=30U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos2 0  _net0 A B _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=30U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net2 Aprime 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos3 0  _net0 B vin _net0 IHP_PDK_nonlinear_components_sg13_lv_pmos w=30U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_pmos4 0  _net1 vin _net3 _net1 IHP_PDK_nonlinear_components_sg13_lv_pmos w=10U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 vin 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=5U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos3 0  vin _net2 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos4 0  Aprime vin 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=15U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

Xsg13_lv_nmos5 0  A HBarre Aprime 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=10U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos6 0  B H _net2 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=12U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
.ENDS
.SUBCKT Diviseur_par_4_symbole _net0 _net1 _net4 

.LIB cornerMOSlv.lib mos_tt


XSUB1 _net2 _net3 INV_2x
XDIVFREQ1 _net3 _net1 _net0 Diviseur_par_2_symbole
XDIVFREQ2 _net4 _net2 _net3 Diviseur_par_2_symbole
.ENDS
.SUBCKT DIV_PAR_256_VF _net12 _net13 V256 

.LIB /home/userproj/microelectronics/PDK/IHP/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt


.LIB cornerMOSlv.lib mos_tt

XSUB2 V4 _net0 Diviseur_par_2_digital_symbole_
V3 _net1 0 DC 1.2
Xsg13_lv_pmos1 0  _net1 _net0 V8 _net1 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  V8 _net0 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
V4 _net2 0 DC 1.2
Xsg13_lv_pmos2 0  _net2 _net3 V16 _net2 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  V16 _net3 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
XSUB4 V16 _net4 Diviseur_par_2_digital_symbole_
V5 _net5 0 DC 1.2
Xsg13_lv_pmos3 0  _net5 _net4 V32 _net5 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos3 0  V32 _net4 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
XSUB5 V32 _net6 Diviseur_par_2_digital_symbole_
V6 _net7 0 DC 1.2
Xsg13_lv_pmos4 0  _net7 _net6 V64 _net7 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos4 0  V64 _net6 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
XSUB6 V64 _net8 Diviseur_par_2_digital_symbole_
V7 _net9 0 DC 1.2
Xsg13_lv_pmos5 0  _net9 _net8 V128 _net9 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos5 0  V128 _net8 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
XSUB7 V128 _net10 Diviseur_par_2_digital_symbole_
V8 _net11 0 DC 1.2
Xsg13_lv_pmos6 0  _net11 _net10 V256 _net11 IHP_PDK_nonlinear_components_sg13_lv_pmos w=2U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos6 0  V256 _net10 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=0.13U ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1


XSUB1 _net13 _net12 V4 Diviseur_par_4_symbole
XSUB8 V8 _net3 Diviseur_par_2_digital_symbole_
.ENDS
.SUBCKT Modele_Inductance _net2 _net1 _net4 
Ls _net0 _net1  2.885N 
Rs _net2 _net0  3.623 tc1=0.0 tc2=0.0 
Csp _net1 _net2  13.69F 
Cox2 _net3 _net1  55.8F 
Rp2 _net4 _net3  18.32 tc1=0.0 tc2=0.0 
Rp1 _net4 _net5  18.32 tc1=0.0 tc2=0.0 
Cox1 _net5 _net2  55.8F 
.ENDS

.SUBCKT IHP_PDK_basic_components_cap_cmim  gnd P1 P2  l=7.0u w=7.0u
X1 P1 P2 cap_cmim l={l} w={w}
.ENDS
  

.SUBCKT IHP_PDK_basic_components_rhigh  gnd P1 P2 w=1.0e-6 l=0.5e-6 m=1
X1 P1 P2 rhigh w={w} l={l} m={m}
.ENDS
  
.SUBCKT symbol _net1 _net3 _net4 VCO= 

.LIB cornerRES.lib res_typ
.LIB cornerCAP.lib cap_typ
.LIB cornerMOSlv.lib mos_tt

XSUB1 _net0 _net1 0 Modele_Inductance
V1 _net0 0 DC 1.2
V6 _net2 0 DC 1.2
Xsg13_lv_nmos4 0  _net5 _net1 _net5 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=200U l=130N ng=20 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos3 0  _net5 _net4 _net5 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=200U l=130N ng=20 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos1 0  _net1 _net4 _net6 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=20U l=130N ng=2 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net4 _net1 _net6 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=20U l=130N ng=2 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos5 0  _net6 _net7 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=10U l=130N ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos6 0  _net7 _net7 0 gnd IHP_PDK_nonlinear_components_sg13_lv_nmos w=1U l=130N ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xcap_cmim2 0  _net4 _net1 IHP_PDK_basic_components_cap_cmim l=18.4U w=18.4U
Xcap_cmim1 0  0 _net7 IHP_PDK_basic_components_cap_cmim l=200U w=200U
Xrhigh1 0  _net2 _net7 IHP_PDK_basic_components_rhigh w=2.1U l=4.1U m=1
Xrhigh2 0  _net3 _net5 IHP_PDK_basic_components_rhigh w=3.1U l=1.6U m=1
XSUB2 _net0 _net4 0 Modele_Inductance

.ENDS

.LIB cornerRES.lib res_typ
.LIB cornerCAP.lib cap_typ
.LIB cornerMOSlv.lib mos_tt

V1 _net0 0 DC 1
XSUB1 _net1 _net2 VOUT DIV_PAR_256_VF
XSUB2 _net2 _net0 _net1 symbol VCO=


.control

tran 5.02513e-10 1e-07 0 
write spice4qucs.tr1.plot v(VOUT)
destroy all
reset

exit
.endc
.END
