* Extracted by KLayout with SG13G2 LVS runset on : 05/06/2025 09:55

.SUBCKT nmos$1
M$1 \$2 \$5 \$3 \$1 sg13_lv_nmos L=0.13u W=100u AS=34p AD=34p PS=200.68u
+ PD=200.68u
.ENDS nmos$1
