*test NETLIST

.SUBCKT TOP
M1 1 2 3 3 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS
