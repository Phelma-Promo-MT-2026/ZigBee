** sch_path: /home/userproj/microelectronics/projects/ZigBee/LVS/xschem/TOP.sch
.subckt TOP

M2 grille grille GND GND sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends
