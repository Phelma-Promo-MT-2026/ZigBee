* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 11:35

.SUBCKT TOP
M$1 \$3 \$4 \$1 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p PS=1.34u
+ PD=0.74u
M$2 \$1 \$4 \$3 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p PS=0.74u
+ PD=1.34u
M$3 \$3 \$4 \$2 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.057p PS=1.28u
+ PD=0.68u
M$4 \$2 \$4 \$3 \$2 sg13_lv_pmos L=0.13u W=0.3u AS=0.057p AD=0.102p PS=0.68u
+ PD=1.28u
.ENDS TOP
