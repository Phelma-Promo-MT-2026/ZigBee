* Extracted by KLayout with SG13G2 LVS runset on : 10/06/2025 11:49

.SUBCKT TOP
M$1 VDD VIN GND GND sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p PS=1.34u
+ PD=1.34u
.ENDS TOP
