* Qucs 25.1.2  /home/userproj/microelectronics/projects/ZigBee/LVS/qucs/cascode/cascode.sch

.SUBCKT IHP_PDK_nonlinear_components_sg13_lv_nmos  gnd d g s b w=0.35u l=0.34u ng=1 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346e-6 z2=0.38e-6 wmin=0.15e-6 rfmode=0 pre_layout=1 mlist=1
X1 d g s b  sg13_lv_nmos w={w} l={l} ng={ng} m={m} as={as} ad={ad} pd={pd} 
+ ps={ps} trise={trise} z1={z1} z2={z2} wmin={wmin} rfmode={rfmode} pre_layout={pre_layout} 
.ENDS
  
.GLOBAL 0:G
Xsg13_lv_nmos1 0  _net0 _net1 _net2 _net2 IHP_PDK_nonlinear_components_sg13_lv_nmos w=100U l=0.130U ng=10 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1
Xsg13_lv_nmos2 0  _net3 _net3 _net0 _net2 IHP_PDK_nonlinear_components_sg13_lv_nmos w=100U l=0.130U ng=10 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1




.END
