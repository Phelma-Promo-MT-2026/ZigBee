* Qucs 25.1.2  /home/userproj/microelectronics/projects/ZigBee/LVS/qucs/nmos_10g_alone/nmos.sch
.GLOBAL 0:G

Xsg13_lv_nmos1 0  Vdd Vin Source 0 IHP_PDK_nonlinear_components_sg13_lv_nmos w=100U l=0.130U ng=10 m=1 as=0 ad=0 pd=0 ps=0 trise=0 z1=0.346E-6 z2=0.38E-6 wmin=0.15E-6 rfmode=0 pre_layout=1

.END
