** sch_path: /home/userproj/microelectronics/projects/ZigBee/LVS/xschem/TOP.sch
**.subckt TOP
XM1 grille grille GND GND sg13_hv_nmos w=1.0u l=0.72u ng=1 m=1 rfmode=1
**.ends
.GLOBAL GND
.end
